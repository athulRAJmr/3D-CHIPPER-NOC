module chipper_tb;
reg [31:0] NORTHIN, SOUTHIN, EASTIN, WESTIN, PEIN,UPIN, DOWNIN;
wire [31:0]NORTHOUT, EASTOUT, SOUTHOUT, WESTOUT, PEOUT, UPOUT, DOWNOUT;
reg inject_request;
wire inject_grant;

chipper #(2'b01, 2'b01,2'b01) Noc_router(NORTHIN, SOUTHIN, EASTIN, WESTIN, UPIN, DOWNIN, PEIN, NORTHOUT, SOUTHOUT, EASTOUT, WESTOUT, UPOUT, DOWNOUT, PEOUT,inject_request, inject_grant);

initial 
begin
  
  #5 NORTHIN <= 32'b01010100111111111111111111111100;
     SOUTHIN <= 32'b11101101111111111111111111111000;
     EASTIN  <= 32'b10100101111111111111111111111000;
     WESTIN  <= 32'b10110000000000000000000000000000;
     UPIN    <= 32'b10110101111111111111111111111000;
     DOWNIN  <= 32'b10110101111111111111111111111000;
     PEIN    <= 32'b01110111111111111111111111111000;
     inject_request <=1'b1;
  
  #5 NORTHIN <= 32'b01000111111111111111111111111000;
     SOUTHIN <= 32'b10101101111111111111111111111000;
     EASTIN  <= 32'b10100101111111111111111111111000;
     WESTIN  <= 32'b11110101111111111111111111111000;
     UPIN    <= 32'b10110101111111111111111111111000;
     DOWNIN  <= 32'b10110101111111111111111111111000;
     PEIN    <= 32'b10110101111111111111111111111000;
     inject_request <=1'b1;
  
  #5 NORTHIN <= 32'b10100101111111111111111111111000;
     SOUTHIN <= 32'b10101101111111111111111111111000;
     EASTIN  <= 32'b10100101111111111111111111111000;
     WESTIN  <= 32'b00110011111111111111111111111000;
     UPIN    <= 32'b10110101111111111111111111111000;
     DOWNIN  <= 32'b10110101111111111111111111111000;
     PEIN    <= 32'b10110101111111111111111111111000;
     inject_request <=1'b1;
  
  #5 NORTHIN <= 32'b10100101111111111111111111111000;
     SOUTHIN <= 32'b10101101111111111111111111111000;
     EASTIN  <= 32'b01010101111111111111111111111000;
     WESTIN  <= 32'b11110101111111111111111111111000;
     UPIN    <= 32'b10110101111111111111111111111000;
     DOWNIN  <= 32'b10110111111111111111111111111000;
     PEIN    <= 32'b10110101111111111111111111111000;
     inject_request <=1'b1;

  

end


initial
begin
 $dumpfile ("chipper.vcd");
 $dumpvars (0, chipper_tb);
$monitor ($time, "NORTHIN =%b, SOUTHIN=%b, EASTIN=%b, WESTIN=%b, PEIN=%b, NORTHOUT=%b, SOUTHOUT=%b, EASTOUT=%b, WESTOUT=%b,PEOUT=%b",
NORTHIN, SOUTHIN, EASTIN, WESTIN, PEIN, NORTHOUT, EASTOUT, SOUTHOUT, WESTOUT, PEOUT );
 #25 $finish;
end
endmodule  